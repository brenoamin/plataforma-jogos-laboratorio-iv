
module sistema_embarcado (
	clk_clk);	

	input		clk_clk;
endmodule
