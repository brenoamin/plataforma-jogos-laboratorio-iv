
module vga (
	clk_clk);	

	input		clk_clk;
endmodule
